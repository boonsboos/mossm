module check

import token
import parse

pub fn check(nodes []parse.Node) {

}