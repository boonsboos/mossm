module parse

