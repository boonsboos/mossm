module parse

import token

pub fn parse(tokens []token.Token) []Node {
	
}