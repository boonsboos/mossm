module parse

pub struct InstructionNode {
	
}

pub struct LabelNode {

}