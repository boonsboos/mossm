module parse

pub type Node = InstructionNode | LabelNode | IdentifierNode

pub struct InstructionNode {
	
}

pub struct LabelNode {

}

pub struct IdentifierNode {

}